module Traffic_light_top(
    input i_clk,                  // Clock input for the entire traffic light system
    input i_reset,                // Asynchronous reset input for initializing or resetting the system
    input i_Vs,                   // Vehicle sensor input to detect vehicles on the side road
    output o_Main_red,            // Output signal for the main road's red light
    output o_Main_yellow,         // Output signal for the main road's yellow light
    output o_Main_green,          // Output signal for the main road's green light
    output o_Side_red,            // Output signal for the side road's red light
    output o_Side_yellow,         // Output signal for the side road's yellow light
    output o_Side_green           // Output signal for the side road's green light
    );

    // Internal signals to connect different modules
    wire [1:0] w_G;               // Gray code output from the sequential logic (current FSM state)
    wire w_Long_trigger;          // Long timer trigger signal from the combinational logic
    wire w_Short_trigger;         // Short timer trigger signal from the combinational logic
    wire w_long_timer;            // Long timer signal generated by the timing circuit
    wire w_short_timer;           // Short timer signal generated by the timing circuit
    wire w_clk;                   // Clock signal used for driving the sequential logic

    // Instantiation of the sequential logic module
    Traffic_Sequential seq_logic (
        .i_Vs(i_Vs),              // Connects the vehicle sensor input to the sequential logic
        .i_clk(w_clk),            // Connects the internal clock to the sequential logic
        .i_Tl(w_long_timer),      // Connects the long timer signal to the sequential logic
        .i_Ts(w_short_timer),     // Connects the short timer signal to the sequential logic
        .i_reset(i_reset),        // Connects the reset signal to the sequential logic
        .o_G(w_G)                 // Outputs the current state as a gray code to the combinational logic
    );

    // Instantiation of the combinational logic module
    Traffic_Combinational comb_logic (
        .i_G(w_G),                // Takes the gray code state from the sequential logic
        .o_Main_red(o_Main_red),  // Controls the main road's red light
        .o_Main_yellow(o_Main_yellow), // Controls the main road's yellow light
        .o_Main_green(o_Main_green),   // Controls the main road's green light
        .o_Side_red(o_Side_red),       // Controls the side road's red light
        .o_Side_yellow(o_Side_yellow), // Controls the side road's yellow light
        .o_Side_green(o_Side_green),   // Controls the side road's green light
        .o_Long_trigger(w_Long_trigger), // Outputs the long timer trigger signal to the timing circuit
        .o_Short_trigger(w_Short_trigger) // Outputs the short timer trigger signal to the timing circuit
    );

    // Instantiation of the timing circuit module
    Traffic_Timing_Circuit timing_circuit (
        .i_clk(i_clk),            // Connects the system clock to the timing circuit
        .i_reset(i_reset),        // Connects the reset signal to the timing circuit
        .i_Long_time(w_Long_trigger),  // Takes the long timer trigger from the combinational logic
        .i_Short_time(w_Short_trigger), // Takes the short timer trigger from the combinational logic
        .o_short_timer(w_short_timer),  // Outputs the short timer signal to the sequential logic
        .o_long_timer(w_long_timer),    // Outputs the long timer signal to the sequential logic
        .o_clk(w_clk)             // Outputs a clock signal that is used by the sequential logic
    );
endmodule

